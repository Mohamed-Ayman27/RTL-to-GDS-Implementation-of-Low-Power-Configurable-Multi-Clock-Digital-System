module CTRL_RX #(
    parameter DATA_WIDTH = 8,
    parameter RF_ADDR    = 4
) (
    input wire CLK,
    input wire RST_
);
    
endmodule